** Profile: "EVM_switching_tb-trans"  [ C:\Users\dwegg\Desktop\Inverter\HW\Simulations\GD_UCC21710\ucc21710-pspicefiles\evm_switching_tb\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ucc21710_trans.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\17.4.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500u 0 10n SKIPBP 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL2= 40
.OPTIONS ITL4= 40
.OPTIONS VNTOL= 1.0m
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\EVM_switching_tb.net" 


.END
